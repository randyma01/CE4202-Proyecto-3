module Modelado (
    input logic [31:0] x,
	 output logic [31:0] y,
	 input logic [31:0] result
);

logic [31:0] a1 = 32'd1;
logic [31:0] b0 = 32'd2;
logic [31:0] b1 = 32'd3;

logic [31:0] w0 = 32'd10; //W inicial
logic [31:0] xmax = 32'd0;//constante -xmax[n]/2

int cont = 0;




    
endmodule
