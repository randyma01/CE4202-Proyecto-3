module Multi (
    input logic [31:0] x,
	 output logic [31:0] y,
	 input logic [31:0] result
);



    
endmodule
