module Modelado (
    
);
    
endmodule