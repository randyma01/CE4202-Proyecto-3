module SumaPF ();

endmodule
