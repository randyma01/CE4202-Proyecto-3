module Modelado (
    input logic [31:0] x,
	 output logic [31:0] y
);

logic a1 = 32'd1;
logic b0 = 32'd2;
logic b1 = 32'd3;

logic w0 = 32'd10;

int cont = 0;

SumaPF sumapf (x[31], x[30:16], x[15:0],x[31], x[30:16], x[15:0])








    
endmodule
